`timescale 1ns / 1ps

module ukladSekwencyjny(
    input clk,
    input start_stop,
    input r, //active 0
    input forw_backw, //active 0
    output reg [3:0] out
  );
  parameter min = 4'b0000;
  parameter max = 4'b1001;
  reg forw_backw_state;
  initial
  begin
    out = max;
    forw_backw_state = 1'b1;  //initially backw
  end

  always @(negedge forw_backw)
  begin
    forw_backw_state = ~ forw_backw_state;
  end
  always@ (posedge clk or negedge r)
  begin
    if(r == 1'b0)
      out = max;
    else if (start_stop == 1'b0)
    begin
      if (forw_backw_state == 1'b0)
      begin
        if(out == max)
          out = min;
        else
          out = out + 1;
      end
      else if (forw_backw_state == 1'b1)
      begin
        if(out == min)
          out = max;
        else
          out = out - 1;
      end
    end
    else
      out=out;
  end
endmodule
